netcdf NDBC46050v3 {
dimensions:
	time = 245448 ;
	bnds = 2 ;
	position = 1 ;
variables:
	float latitude ;
		latitude:units = "degrees_north" ;
		latitude:long_name = "latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:valid_min = 44.656 ;
		latitude:valid_max = 44.656 ;
		latitude:axis = "Y" ;
	float longitude(position) ;
		longitude:units = "degrees_east" ;
		longitude:long_name = "longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:valid_min = 235.474 ;
		longitude:valid_max = 235.474 ;
		longitude:axis = "X" ;
	float time(time) ;
		time:units = "hours since 1970-01-01" ;
		time:calendar = "gregorian" ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
		time:valid_min = 149016. ;
		time:valid_max = 394463. ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
	float depth(position) ;
		depth:units = "meters" ;
		depth:long_name = "Depth of each measurement" ;
		depth:standard_name = "depth" ;
		depth:valid_min = -1. ;
		depth:valid_max = -1. ;
		depth:axis = "Z" ;
		depth:positive = "up" ;
	int station_name(position) ;
		station_name:long_name = "station name" ;
		station_name:cf_role = "timeseries_id" ;
		station_name:units = "1" ;
	float time_bnds(time, bnds) ;
		time_bnds:units = "hours since 1970-01-01" ;
		time_bnds:long_name = "time cell boundaries" ;
	float sea_water_temperature(time) ;
		sea_water_temperature:_FillValue = -9999.f ;
		sea_water_temperature:units = "degree_Celsius" ;
		sea_water_temperature:cell_methods = "time: mean (interval: 1 hour comment: time indicates center hour)" ;
		sea_water_temperature:long_name = "Hourly Sea Water Temperature" ;
		sea_water_temperature:standard_name = "sea_water_temperature" ;
		sea_water_temperature:coordinates = "longitude latitude time depth" ;
		sea_water_temperature:sensor_mount = "mounted on mooring bridal" ;
		sea_water_temperature:valid_min = -2. ;
		sea_water_temperature:valid_max = 30. ;

// global attributes:
		:title = "Hourly NDBC 46050 data" ;
		:publisher_name = "Craig Risien" ;
		:publisher_email = "crisien@coas.oregonstate.edu" ;
		:institution = "Oregon State University, College of Earth, Ocean, and Atmospheric Sciences" ;
		:date_created = "2015-11-13T12:51:22" ;
		:date_modified = "2015-11-13T12:51:22" ;
		:history = "Quality controlled at NOAA NDBC" ;
		:time_coverage_start = "1987-01-01T00:00:00" ;
		:time_coverage_end = "2014-12-31T23:00:00" ;
		:time_coverage_resolution = "hourly averages" ;
		:geospatial_lat_min = 44.656 ;
		:geospatial_lat_max = 44.656 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_min = 235.474 ;
		:geospatial_lon_max = 235.474 ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_vertical_min = -1. ;
		:geospatial_vertical_max = -1. ;
		:geospatial_vertical_units = "meters" ;
		:geospatial_vertical_resolution = "point" ;
		:geospatial_vertical_positive = "up" ;
		:keywords = "sea surface temperature, ndbc, noaa" ;
		:keyword_vocabulary = "GCMD" ;
		:Conventions = "CF-1.6" ;
		:comments = "no comment" ;
		:cdm_data_type = "Station" ;
		:featureType = "timeSeries" ;
		:data_type = "NDBC time-series data" ;
		:area = "North Pacific Ocean" ;
		:license = "Follows NDBC standards. Data available free of charge. User assumes all risk for use of data. User must display citation in any publication or product using data." ;
		:citation = "These data were collected and made freely available by NOAA NDBC" ;
		:acknowledgement = "These data were collected and made freely available by NOAA NDBC" ;
		:wmo_platform_code = "46050" ;
		:summary = "Quality controlled NDBC Station data that have been repackaged and distributed by NANOOS" ;
		:naming_authority = "NOAA NDBC" ;
}
