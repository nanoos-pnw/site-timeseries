netcdf NDBC46029 {
dimensions:
	time = 280512 ;
	bnds = 2 ;
variables:
	float latitude ;
		latitude:units = "degrees_north" ;
		latitude:long_name = "latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:valid_min = 46.159 ;
		latitude:valid_max = 46.159 ;
		latitude:axis = "Y" ;
	float longitude ;
		longitude:units = "degrees_east" ;
		longitude:long_name = "longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:valid_min = 235.486 ;
		longitude:valid_max = 235.486 ;
		longitude:axis = "X" ;
	float time(time) ;
		time:units = "hours since 1970-01-01" ;
		time:calendar = "gregorian" ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
		time:valid_min = 122712. ;
		time:valid_max = 403223. ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
	float depth_sst ;
		depth_sst:units = "meters" ;
		depth_sst:long_name = "Depth of SST measurements" ;
		depth_sst:standard_name = "depth" ;
		depth_sst:valid_min = -0.6 ;
		depth_sst:valid_max = -0.6 ;
		depth_sst:axis = "Z" ;
		depth_sst:positive = "up" ;
	float depth_atmp ;
		depth_atmp:units = "meters" ;
		depth_atmp:long_name = "Height of air temperature measurements" ;
		depth_atmp:standard_name = "depth" ;
		depth_atmp:valid_min = 4. ;
		depth_atmp:valid_max = 4. ;
		depth_atmp:axis = "Z" ;
		depth_atmp:positive = "up" ;
	float depth_wnd ;
		depth_wnd:units = "meters" ;
		depth_wnd:long_name = "Height of wind measurements" ;
		depth_wnd:standard_name = "depth" ;
		depth_wnd:valid_min = 5. ;
		depth_wnd:valid_max = 5. ;
		depth_wnd:axis = "Z" ;
		depth_wnd:positive = "up" ;
	float depth_press ;
		depth_press:units = "meters" ;
		depth_press:long_name = "Height of barometric pressure measurements" ;
		depth_press:standard_name = "depth" ;
		depth_press:valid_min = 0. ;
		depth_press:valid_max = 0. ;
		depth_press:axis = "Z" ;
		depth_press:positive = "up" ;
	float depth_wav ;
		depth_wav:units = "meters" ;
		depth_wav:long_name = "Height of wave measurements" ;
		depth_wav:standard_name = "depth" ;
		depth_wav:valid_min = 0. ;
		depth_wav:valid_max = 0. ;
		depth_wav:axis = "Z" ;
		depth_wav:positive = "up" ;
	int station_name ;
		station_name:long_name = "station name" ;
		station_name:cf_role = "timeseries_id" ;
		station_name:units = "1" ;
	float time_bnds(time, bnds) ;
		time_bnds:units = "hours since 1970-01-01" ;
		time_bnds:long_name = "time cell boundaries" ;
		time_bnds:calendar = "gregorian" ;
	float sea_water_temperature(time) ;
		sea_water_temperature:_FillValue = -9999.f ;
		sea_water_temperature:units = "K" ;
		sea_water_temperature:cell_methods = "time: mean (interval: 1 hour comment: time indicates center hour)" ;
		sea_water_temperature:long_name = "Hourly Sea Water Temperature" ;
		sea_water_temperature:standard_name = "sea_water_temperature" ;
		sea_water_temperature:coordinates = "longitude latitude time depth_sst" ;
		sea_water_temperature:sensor_mount = "mounted on mooring bridal" ;
		sea_water_temperature:valid_min = 271.15 ;
		sea_water_temperature:valid_max = 303.15 ;
	float air_temperature(time) ;
		air_temperature:_FillValue = -9999.f ;
		air_temperature:units = "K" ;
		air_temperature:cell_methods = "time: mean (interval: 1 hour comment: time indicates center hour)" ;
		air_temperature:long_name = "Hourly Air Temperature" ;
		air_temperature:standard_name = "air_temperature" ;
		air_temperature:coordinates = "longitude latitude time depth_atmp" ;
		air_temperature:sensor_mount = "mounted on the buoy tower" ;
		air_temperature:valid_min = 243.15 ;
		air_temperature:valid_max = 303.15 ;
	float air_pressure(time) ;
		air_pressure:_FillValue = -9999.f ;
		air_pressure:units = "Pa" ;
		air_pressure:cell_methods = "time: mean (interval: 1 hour comment: time indicates center hour)" ;
		air_pressure:long_name = "Hourly Air Pressure" ;
		air_pressure:standard_name = "air_pressure_at_sea_level" ;
		air_pressure:coordinates = "longitude latitude time depth_press" ;
		air_pressure:sensor_mount = "mounted on the buoy tower" ;
		air_pressure:valid_min = 95000. ;
		air_pressure:valid_max = 105000. ;
	float wind_speed(time) ;
		wind_speed:_FillValue = -9999.f ;
		wind_speed:units = "m s-1" ;
		wind_speed:cell_methods = "time: mean (interval: 1 hour comment: time indicates center hour)" ;
		wind_speed:long_name = "Hourly Wind Speed" ;
		wind_speed:standard_name = "wind_speed" ;
		wind_speed:coordinates = "longitude latitude time depth_wnd" ;
		wind_speed:sensor_mount = "mounted on the buoy tower" ;
		wind_speed:valid_min = 0. ;
		wind_speed:valid_max = 60. ;
	float wind_speed_gust(time) ;
		wind_speed_gust:_FillValue = -9999.f ;
		wind_speed_gust:units = "m s-1" ;
		wind_speed_gust:cell_methods = "time: mean (interval: 1 hour comment: time indicates center hour)" ;
		wind_speed_gust:long_name = "Hourly Wind Speed Gust" ;
		wind_speed_gust:standard_name = "wind_speed_of_gust" ;
		wind_speed_gust:coordinates = "longitude latitude time depth_wnd" ;
		wind_speed_gust:sensor_mount = "mounted on the buoy tower" ;
		wind_speed_gust:valid_min = 0. ;
		wind_speed_gust:valid_max = 60. ;
	float wind_direction(time) ;
		wind_direction:_FillValue = -9999.f ;
		wind_direction:units = "degree" ;
		wind_direction:cell_methods = "time: mean (interval: 1 hour comment: time indicates center hour)" ;
		wind_direction:long_name = "Hourly Wind Direction" ;
		wind_direction:standard_name = "wind_from_direction" ;
		wind_direction:coordinates = "longitude latitude time depth_wnd" ;
		wind_direction:sensor_mount = "mounted on the buoy tower" ;
		wind_direction:valid_min = 0. ;
		wind_direction:valid_max = 360. ;
	float significant_wave_height(time) ;
		significant_wave_height:_FillValue = -9999.f ;
		significant_wave_height:units = "m" ;
		significant_wave_height:cell_methods = "time: mean (interval: 1 hour comment: time indicates center hour)" ;
		significant_wave_height:long_name = "Hourly Significant Height of Wind and Swell Waves" ;
		significant_wave_height:standard_name = "sea_surface_wave_significant_height" ;
		significant_wave_height:coordinates = "longitude latitude time depth_wav" ;
		significant_wave_height:sensor_mount = "mounted in the buoy" ;
		significant_wave_height:valid_min = 0. ;
		significant_wave_height:valid_max = 20. ;
	float average_wave_period(time) ;
		average_wave_period:_FillValue = -9999.f ;
		average_wave_period:units = "s" ;
		average_wave_period:cell_methods = "time: mean (interval: 1 hour comment: time indicates center hour)" ;
		average_wave_period:long_name = "Hourly Average Wave Period" ;
		average_wave_period:standard_name = "average_wave_period" ;
		average_wave_period:coordinates = "longitude latitude time depth_wav" ;
		average_wave_period:sensor_mount = "mounted in the buoy" ;
		average_wave_period:valid_min = 0. ;
		average_wave_period:valid_max = 30. ;
	float dominant_wave_period(time) ;
		dominant_wave_period:_FillValue = -9999.f ;
		dominant_wave_period:units = "s" ;
		dominant_wave_period:cell_methods = "time: mean (interval: 1 hour comment: time indicates center hour)" ;
		dominant_wave_period:long_name = "Hourly Dominant Wave Period" ;
		dominant_wave_period:standard_name = "dominant_wave_period" ;
		dominant_wave_period:coordinates = "longitude latitude time depth_wav" ;
		dominant_wave_period:sensor_mount = "mounted in the buoy" ;
		dominant_wave_period:valid_min = 0. ;
		dominant_wave_period:valid_max = 30. ;
	float mean_wave_direction(time) ;
		mean_wave_direction:_FillValue = -9999.f ;
		mean_wave_direction:units = "degree" ;
		mean_wave_direction:cell_methods = "time: mean (interval: 1 hour comment: time indicates center hour)" ;
		mean_wave_direction:long_name = "Hourly Mean Wave Direction" ;
		mean_wave_direction:standard_name = "sea_surface_wave_from_direction" ;
		mean_wave_direction:coordinates = "longitude latitude time depth_wav" ;
		mean_wave_direction:sensor_mount = "mounted in the buoy" ;
		mean_wave_direction:valid_min = 0. ;
		mean_wave_direction:valid_max = 360. ;

// global attributes:
		:title = "Hourly NDBC 46029 data" ;
		:publisher_name = "Craig Risien" ;
		:publisher_email = "crisien@coas.oregonstate.edu" ;
		:institution = "Oregon State University, College of Earth, Ocean, and Atmospheric Sciences" ;
		:date_created = "2015-11-17T12:58:28" ;
		:date_modified = "2015-11-17T12:58:28" ;
		:history = "Quality controlled at NOAA NDBC" ;
		:time_coverage_start = "1984-01-01T00:00:00" ;
		:time_coverage_end = "2015-12-31T23:00:00" ;
		:time_coverage_resolution = "hourly averages" ;
		:geospatial_lat_min = 46.159 ;
		:geospatial_lat_max = 46.159 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_min = 235.486 ;
		:geospatial_lon_max = 235.486 ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_vertical_min = -0.6 ;
		:geospatial_vertical_max = 5. ;
		:geospatial_vertical_units = "meters" ;
		:geospatial_vertical_resolution = "point" ;
		:geospatial_vertical_positive = "up" ;
		:keywords = "ndbc, noaa, nanoos, sea surface temperature, wind speed, wind direction, wave height, wave period, wave direction, air temperature, barometric pressure" ;
		:keyword_vocabulary = "GCMD" ;
		:Conventions = "CF-1.6" ;
		:comments = "no comment" ;
		:cdm_data_type = "Station" ;
		:featureType = "timeSeries" ;
		:data_type = "NDBC time-series data" ;
		:area = "North Pacific Ocean" ;
		:license = "Follows NDBC standards. Data available free of charge. User assumes all risk for use of data. User must display citation in any publication or product using data." ;
		:citation = "These data were collected and made freely available by NOAA NDBC" ;
		:acknowledgement = "These data were collected and made freely available by NOAA NDBC" ;
		:wmo_platform_code = "46029" ;
		:summary = "Quality controlled NDBC Station data that have been repackaged and distributed by NANOOS" ;
		:naming_authority = "NOAA NDBC" ;
}
