netcdf OS_PAP-3_201205_P_deepTS {
dimensions:
	TIME = 16767 ;
	DEPTH = 1 ;
	LATITUDE = 1 ;
	LONGITUDE = 1 ;
variables:
	double TIME(TIME) ;
		TIME:description = "Date and Time from Matlab" ;
		TIME:long_name = "time" ;
		TIME:standard_name = "time" ;
		TIME:units = "days since 1950-01-01T00:00:00Z" ;
		TIME:conventions = "Relative julian days with decimal part (as parts of the day)" ;
		TIME:valid_min = 0. ;
		TIME:valid_max = 90000. ;
		TIME:QC_indicator = "good_data" ;
		TIME:processing_level = "Instrument data that has been converted to geophysical values" ;
		TIME:uncertainty = 5.e-06 ;
		TIME:axis = "T" ;
	float DEPTH(DEPTH) ;
		DEPTH:long_name = "Depth of each measurement" ;
		DEPTH:standard_name = "depth" ;
		DEPTH:units = "meters" ;
		DEPTH:positive = "down" ;
		DEPTH:valid_min = 0. ;
		DEPTH:valid_max = 12000. ;
		DEPTH:comment = "These are nominal values. Use PRES to derive time-varying depths of instruments, as the mooring may tilt in ambient currents." ;
		DEPTH:QC_indicator = "good_data" ;
		DEPTH:processing_level = "Instrument data that has been converted to geophysical values" ;
		DEPTH:uncertainty = "0" ;
		DEPTH:axis = "Z" ;
		DEPTH:reference = "WGS84" ;
		DEPTH:coordinate_reference_frame = "urn:ogc:def:crs:EPSG::4326" ;
	float LATITUDE(LATITUDE) ;
		LATITUDE:QC_indicator = "good_data" ;
		LATITUDE:processing_level = "Instrument data that has been converted to geophysical values" ;
		LATITUDE:long_name = "Latitude of each location" ;
		LATITUDE:standard_name = "latitude" ;
		LATITUDE:units = "degrees_north" ;
		LATITUDE:valid_min = -90. ;
		LATITUDE:valid_max = 90. ;
		LATITUDE:comment = "LATITUDE Latitude for each point" ;
		LATITUDE:ancillary_variables = "LATITUDE_QC" ;
		LATITUDE:uncertainty = 0.05 ;
		LATITUDE:axis = "Y" ;
	float LONGITUDE(LONGITUDE) ;
		LONGITUDE:QC_indicator = "good_data" ;
		LONGITUDE:procedding_level = "Instrument data that has been converted to geophysical values" ;
		LONGITUDE:long_name = "Longitude of each location" ;
		LONGITUDE:standard_name = "longitude" ;
		LONGITUDE:units = "degrees_east" ;
		LONGITUDE:valid_min = -180. ;
		LONGITUDE:valid_max = 180. ;
		LONGITUDE:comment = "LONGITUDE Longitude for each point" ;
		LONGITUDE:ancillary_variables = "LONGITUDE_QC" ;
		LONGITUDE:uncertainty = 0.05 ;
		LONGITUDE:axis = "X" ;
	float TEMP(TIME, DEPTH) ;
		TEMP:long_name = "Temperature" ;
		TEMP:standard_name = "sea_water_temperature" ;
		TEMP:valid_min = 2. ;
		TEMP:valid_max = 100. ;
		TEMP:comment = "Temperature in Degrees Celsius at nominal depths of 4850 meter(s)" ;
		TEMP:units = "degree_Celsius" ;
		TEMP:coordinates = "TIME DEPTH LATITUDE LONGITUDE" ;
		TEMP:sensor_depth = "4850  m(s)" ;
		TEMP:sensor_mount = "mounted on mooring line" ;
		TEMP:sensor_orientation = "vertical" ;
		TEMP:_FillValue = 99999.f ;
		TEMP:DM_indicator = "P" ;
		TEMP:sensor_name = "Seabird:Seabird SBE 37-IMP with pressure sensor; with Pump  " ;
		TEMP:sensor_serial_number = "9477, " ;
		TEMP:accuracy = 0.003 ;
		TEMP:resolution = 0.001 ;
		TEMP:cell_methods = "TIME: point DEPTH: point" ;
		TEMP:ancillary_variables = "TEMP_QC PRES" ;
		TEMP:processing_level = "Instrument data that has been converted to geophysical values" ;
	byte TEMP_QC(TIME, DEPTH) ;
		TEMP_QC:name = "TEMP_QC" ;
		TEMP_QC:long_name = "quality flag for Temperature in Degrees Celsius at nominal depths of 4850 meter(s)" ;
		TEMP_QC:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		TEMP_QC:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used nominal_value interpolated_value missing_value" ;
		TEMP_QC:coordinates = "TIME DEPTH LATITUDE LONGITUDE" ;
	float CNDC(TIME, DEPTH) ;
		CNDC:long_name = "sea water electrical conductivity" ;
		CNDC:standard_name = "sea_water_electrical_conductivity" ;
		CNDC:valid_min = 25. ;
		CNDC:valid_max = 45. ;
		CNDC:comment = "Conductivity in mS/cm at nominal depths of 4850 meter(s)" ;
		CNDC:units = "mS/cm" ;
		CNDC:coordinates = "TIME DEPTH LATITUDE LONGITUDE" ;
		CNDC:sensor_depth = "4850  m(s)" ;
		CNDC:sensor_mount = "mounted on mooring line" ;
		CNDC:sensor_orientation = "vertical" ;
		CNDC:_FillValue = 99999.f ;
		CNDC:DM_indicator = "P" ;
		CNDC:sensor_name = "Seabird:Seabird SBE 37-IMP with pressure sensor; with Pump  " ;
		CNDC:sensor_serial_number = "9477, " ;
		CNDC:accuracy = 0.02 ;
		CNDC:resolution = 0.001 ;
		CNDC:cell_methods = "TIME: point DEPTH: point" ;
		CNDC:ancillary_variables = "CNDC_QC PRES" ;
		CNDC:processing_level = "Instrument data that has been converted to geophysical values" ;
	byte CNDC_QC(TIME, DEPTH) ;
		CNDC_QC:name = "CNDC_QC" ;
		CNDC_QC:long_name = "quality flag for Conductivity in mS/cm at nominal depths of 4850 meter(s)" ;
		CNDC_QC:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		CNDC_QC:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used nominal_value interpolated_value missing_value" ;
		CNDC_QC:coordinates = "TIME DEPTH LATITUDE LONGITUDE" ;
	float PSAL(TIME, DEPTH) ;
		PSAL:long_name = "sea water salinity" ;
		PSAL:standard_name = "sea_water_practical_salinity" ;
		PSAL:valid_min = 29. ;
		PSAL:valid_max = 40. ;
		PSAL:comment = "Practical PSAL Units for each nominal depth(s) of 4850 meter(s)" ;
		PSAL:units = "1" ;
		PSAL:coordinates = "TIME DEPTH LATITUDE LONGITUDE" ;
		PSAL:sensor_depth = "4850  m(s)" ;
		PSAL:sensor_mount = "mounted on mooring line" ;
		PSAL:sensor_orientation = "vertical" ;
		PSAL:_FillValue = 99999.f ;
		PSAL:DM_indicator = "P" ;
		PSAL:sensor_name = "Seabird:Seabird SBE 37-IMP with pressure sensor; with Pump  " ;
		PSAL:sensor_serial_number = "9477, " ;
		PSAL:accuracy = 0.25 ;
		PSAL:resolution = 0.03 ;
		PSAL:cell_methods = "TIME: point DEPTH: point" ;
		PSAL:ancillary_variables = "PSAL_QC PRES" ;
		PSAL:processing_level = "Instrument data that has been converted to geophysical values" ;
	byte PSAL_QC(TIME, DEPTH) ;
		PSAL_QC:name = "PSAL_QC" ;
		PSAL_QC:long_name = "quality flag for Practical PSAL Units for each nominal depth(s) of 4850 meter(s)" ;
		PSAL_QC:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		PSAL_QC:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used nominal_value interpolated_value missing_value" ;
		PSAL_QC:coordinates = "TIME DEPTH LATITUDE LONGITUDE" ;
	float PRES(TIME, DEPTH) ;
		PRES:long_name = "sea_water_pressure" ;
		PRES:standard_name = "sea_water_pressure" ;
		PRES:valid_min = 0. ;
		PRES:valid_max = 6000. ;
		PRES:comment = "PRES (dbar) at nominal depths of 4850 meter(s)" ;
		PRES:units = "decibar" ;
		PRES:coordinates = "TIME DEPTH LATITUDE LONGITUDE" ;
		PRES:sensor_depth = "4850  m(s)" ;
		PRES:sensor_mount = "mounted on mooring line" ;
		PRES:sensor_orientation = "vertical" ;
		PRES:_FillValue = 99999.f ;
		PRES:DM_indicator = "P" ;
		PRES:sensor_name = "Seabird:Seabird SBE 37-IMP with pressure sensor; with Pump  " ;
		PRES:sensor_serial_number = "9477, " ;
		PRES:accuracy = 0.25 ;
		PRES:resolution = 0.03 ;
		PRES:cell_methods = "TIME: point DEPTH: point" ;
		PRES:ancillary_variables = "PRES_QC" ;
		PRES:processing_level = "Instrument data that has been converted to geophysical values" ;
	byte PRES_QC(TIME, DEPTH) ;
		PRES_QC:name = "PRES_QC" ;
		PRES_QC:long_name = "quality flag for PRES (dbar) at nominal depths of 4850 meter(s)" ;
		PRES_QC:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		PRES_QC:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used nominal_value interpolated_value missing_value" ;
		PRES_QC:coordinates = "TIME DEPTH LATITUDE LONGITUDE" ;

// global attributes:
		:summary = "FixO3 Fixed-point Open Ocean ObservatoriesEU Framework 7 programme (FP7/2007-2013) grant agreement No.312463" ;
		:site_code = "PAP" ;
		:platform_code = "PAP-3" ;
		:data_mode = "P" ;
		:title = "OceanSITES PAP in-situ data" ;
		:naming_authority = "OceanSITES" ;
		:id = "OS_PAP-3_201205_P_deepTS" ;
		:name = "OS_PAP-3_201205_P_deepTS" ;
		:wmo_platform_code = "62442" ;
		:source = "Mooring observation" ;
		:principal_investigator = "Richard Lampitt" ;
		:principal_investigator_email = "R.Lampitt@noc.ac.uk" ;
		:principal_investigator_url = "https://noc.ac.uk/people/rsl" ;
		:institution = "NOC" ;
		:project = "FixO3" ;
		:array = "PAP-SO" ;
		:network = "FixO3" ;
		:keywords_vocabulary = "SeaDataNet Parameter Discovery Vocabulary" ;
		:keywords = "WC_Temp, WC_Sal,http://vocab.nerc.ac.uk/collection/P02/current/TEMP/,http://vocab.nerc.ac.uk/collection/P02/current/PSAL/" ;
		:comment = "no comment" ;
		:area = "North Atlantic Ocean" ;
		:geospatial_lat_min = "48" ;
		:geospatial_lat_max = "50" ;
		:geospatial_lat_units = "degree_north" ;
		:geospatial_lon_min = "-16" ;
		:geospatial_lon_max = "-17" ;
		:geospatial_lon_units = "degree_east" ;
		:geospatial_vertical_min = "4850" ;
		:geospatial_vertical_max = "4850" ;
		:geospatial_vertical_positive = "down" ;
		:geospatial_vertical_units = "meter" ;
		:time_coverage_start = "2012-05-05T12:00:01Z" ;
		:time_coverage_end = "2013-04-19T19:00:01Z" ;
		:time_coverage_duration = "P349D" ;
		:time_coverage_resolution = "PT30M" ;
		:cdm_data_type = "Station" ;
		:featureType = "timeSeries" ;
		:data_type = "OceanSITES time-series data" ;
		:format_version = "1.3" ;
		:Conventions = "CF-1.6" ;
		:netcdf_version = "3.5" ;
		:publisher_name = "Maureen Pagnani" ;
		:publisher_email = "m.pagnani at bodc.ac.uk" ;
		:publisher_url = "http://www.fixo3.eu" ;
		:references = " http://www.fixo3.eu, http://www.oceansites.org, http://www.coriolis.eu.org, http://www.eurosites.info" ;
		:institution_references = " http://noc.ac.uk" ;
		:data_assembly_center = "FixO3 DAC" ;
		:update_interval = "void" ;
		:license = "Follows CLIVAR (Climate Varibility and Predictability) standards, cf. http://www.clivar.org/data/data_policy.php. Data available free of charge. User assumes all risk for use of data. User must display citation in any publication or product using data. User must contact PI prior to any commercial use of data." ;
		:citation = "These data were collected and made freely available from the Porcupine Abyssal Plain (PAP) Observatory and the UK national programs that contribute to it, together with European Projects (FixO3, EuroSITES, MERSEA, ANIMATE) that have supported it, and the OceanSITES project." ;
		:acknowledgement = "These data were collected and made freely available from the Porcupine Abyssal Plain (PAP) Observatory and the UK national programs that contribute to it, together with European Projects (FixO3, EuroSITES, MERSEA, ANIMATE) that have supported it, and the OceanSITES project." ;
		:date_created = "2015-06-04T17:25:53Z" ;
		:date_modified = "2015-06-04T17:25:53Z" ;
		:history = "Near real-time processed quality controlled at DAC" ;
		:processing_level = "Instrument data that has been converted to geophysical values" ;
		:QC_indicator = "1" ;
		:contributor_name = "Corinne Pebody" ;
		:contributor_role = "Editor" ;
		:contributor_email = "cawo@noc.ac.uk" ;
}
